module prac_tb();
	reg [255:0] p, q;

	wire [232:0] result;
		ks256 dut(.p(p),.q(q),.result(result));
	initial 
		begin
			$monitor($time,"P = %b, Q = %b, Y = %b",p,q,result);
			#5 p = 256'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111;
			#5 q = 256'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
			#5 $finish;
		end
endmodule


